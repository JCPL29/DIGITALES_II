library verilog;
use verilog.vl_types.all;
entity outputports_vlg_vec_tst is
end outputports_vlg_vec_tst;
