library verilog;
use verilog.vl_types.all;
entity ALUtest_vlg_vec_tst is
end ALUtest_vlg_vec_tst;
